module Exercise1(input A, output x, output y);
    assign x = A;
	 assign y = !A;
endmodule
