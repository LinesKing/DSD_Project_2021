`include "CPU.vh"

// // Step 2 of Stage 5:
// // 	Asynchronous ROM (Program Memory)
//module AsyncROM(input [7:0] addr, output reg [34:0] data);
//	always @(addr)
//		case (addr)
//			0: data = {`MOV, `PUR, `NUM, 8'd 1, `REG, `DOUT, `N8};
//			1: data = {`MOV, `PUR, `NUM, 8'd 3, `REG, `DOUT, `N8};
//			2: data = {`MOV, `PUR, `NUM, 8'd 5, `REG, `DOUT, `N8};
//			3: data = {`MOV, `PUR, `NUM, 8'd 7, `REG, `DOUT, `N8};
//			4: data = {`MOV, `PUR, `NUM, 8'd 9, `REG, `DOUT, `N8};
//			5: data = {`MOV, `PUR, `NUM, 8'd 11, `REG, `DOUT, `N8};
//			6: data = {`MOV, `PUR, `NUM, 8'd 13, `REG, `DOUT, `N8};
//			7: data = {`MOV, `PUR, `NUM, 8'd 15, `REG, `DOUT, `N8};
//			8: data = {`MOV, `PUR, `NUM, 8'd 17, `REG, `DOUT, `N8};
//			9: data = {`MOV, `PUR, `NUM, 8'd 19, `REG, `DOUT, `N8};
//			default: data = 35'b0; // Default instruction is a NOP
//		endcase
//endmodule

module AsyncROM(input [7:0] addr, output reg [34:0] data);
	always @(addr)
		case (addr)
			0: data = set(`DOUT, 1);
			4: data = acc(`SMT, `DOUT, -2);
			8: data = atc(`OFLW, 16);
			12: data = jmp(4);
			16: data = set(`DOUT, 250);
			20: data = acc(`UAD, `DOUT, 1);
			24: data = atc(`OFLW, 8);
			28: data = jmp(20);
			default: data = 35'b0; // NOP
			1, 5, 9, 13, 17, 21, 25: data = mov(`FLAG, `GOUT);
		endcase
		
	function [34:0] set;
		input [7:0] reg_num;
		input [7:0] value;
		set = {`MOV, `PUR, `NUM, value, `REG, reg_num, `N8};
	endfunction
	
	function [34:0] mov;
		input [7:0] src_reg;
		input [7:0] dst_reg;
		mov = {`MOV, `PUR, `REG, src_reg, `REG, dst_reg, `N8};
	endfunction
	
	function [34:0] jmp;
		input [7:0] addr;
		jmp = {`JMP, `UNC, `N10, `N10, addr};
	endfunction
	
	function [34:0] atc;
		input [2:0] bit;
		input [7:0] addr;
		atc = {`ATC, bit, `N10, `N10, addr};
	endfunction
	
	function [34:0] acc;
		input [2:0] op;
		input [7:0] reg_num;
		input [7:0] value;
		acc = {`ACC, op, `REG, reg_num, `NUM, value, `N8};
	endfunction
	
	// Stage 11: Setting and Clearing Individual Bits
	function [34:0] set_bit;
		input [7:0] reg_num;
		input [2:0] bit;
		set_bit = {`ACC, `OR, `REG, reg_num, `NUM, 8'b1 << bit, `N8};
	endfunction
	
	function [34:0] clr_bit;
		input [7:0] reg_num;
		input [2:0] bit;
		clr_bit = {`ACC, `AND, `REG, reg_num, `NUM, ~(8'b1 << bit), `N8};
	endfunction

endmodule
